* TLC27L2 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 07/10/90 AT 15:01
* REV (N/A)      SUPPLY VOLTAGE: 5V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TLC27L2  1 2 3 4 5
*
  C1   11 12 10.12E-12
  C2    6  7 15.00E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  FB 7 99 POLY(5) VB VC VE VLP VLN 0 419.1E6 -70E6 70E6 70E6 -70E6
  GA    6  0 11 12 7.069E-6
  GCM 0  6 10 99 282.0E-12
  HLIM 90  0 VLIM 1K
  ISS   3 10 DC 450.0E-9
  J1   11  2 10 JX
  J2   12  1 10 JX
  R2    6  9 100.0E3
  RD1 60 11 141.5E3
  RD2 60 12 141.5E3
  RO1   8  5 85
  RO2   7 99 85
  RP  3 4 523.6E3
  RSS  10 99 444.4E6
  VAD  60 4 -.5
  VB    9  0 DC 0
  VC 3 53 DC 1.470
  VE   54  4 DC .57
  VLIM  7  8 DC 0
  VLP  91  0 DC 20
  VLN   0 92 DC 20
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=300.0E-15 BETA=222.1E-6 VTO=.027)
.ENDS
