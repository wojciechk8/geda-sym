*
*******************************************
*
*BZX84-C5V1
*
*NXP Semiconductors
*
*Voltage regulator diode
*
*
*
*
*
*VFmax = 0,9V @ IF = 10mA
*IRmax = 2�A  @ VR = 2V
*
*VZmax = 5,4V @ IZ = 5mA
*
*
*
*Ptot  = 250mW
*
*
*
*Package pinning does not match Spice model pinning.
*Package: SOT23 (TO236AB)
*
*Package Pin 1: Anode
*Package Pin 2: not connected
*Package Pin 3: Cathode
*
*
*Extraction date (week/year): 01/2016
*Simulator: SPICE2
*
*******************************************
*
.SUBCKT BZX84_C5V1 1 2
 R1 1 2 1E+011
 D1 1 2
 + DIODE1
 D2 3 1
 + DIODE2
 VZ 2 3 0.1
*
*The resistor R1, the diode D2 and
*VZ do not reflect
*physical devices but improve
*only modeling in the reverse
*mode of operation.
*
 .MODEL DIODE1 D
 + IS = 1E-014
 + N = 1.1
 + BV = 4.8
 + IBV = 1E-009
 + RS = 0.2
 + CJO = 1.2E-010
 + VJ = 0.6
 + M = 0.31
 + FC = 0.5
 + TT = 0
 + EG = 1.1
 + XTI = 3
 .MODEL DIODE2 D
 + IS = 3E-011
 + N = 9.5
 + RS = 30
 .ENDS
*
