*---------- DMC2400UV Spice Model ----------

*NMOS
.SUBCKT DMC2400UV_NMOS 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3  NMOS  L = 1E-006  W = 1E-006 
RD 10 1 0.1925 
RS 30 3 0.001 
RG 20 2 68 
CGS 2 3 3.272E-011 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1  VFB 1 
CGD 13 14 6.7E-011 
R1 13 0 1 
D1 12 13  DLIM 
DDG 15 14  DCGD 
R2 12 15 1 
D2 15 0  DLIM 
DSD 3 10  DSUB 
.MODEL NMOS NMOS  LEVEL = 3  VMAX = 1E+006  ETA = 0.01  VTO = 0.9058 
+ TOX = 6E-008  NSUB = 1E+016  KP = 3.223  U0 = 400  KAPPA = 15.35 
.MODEL DCGD D  CJO = 1.94E-011  VJ = 0.1108  M = 0.3101 
.MODEL DSUB D  IS = 1E-009  N = 1.905  RS = 0.02633  BV = 25  CJO = 5.066E-012  VJ = 0.1753  M = 0.2672 
.MODEL DLIM D  IS = 0.0001 
.ENDS


*PMOS
.SUBCKT DMC2400UV_PMOS 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3  PMOS  L = 1E-006  W = 1E-006 
RD 10 1 0.4041 
RS 30 3 0.001 
RG 20 2 14.3 
CGS 2 3 4.178E-011 
EGD 12 30 2 1 1 
VFB 14 30 0 
FFB 2 1  VFB 1 
CGD 13 14 5.7E-011 
R1 13 30 1 
D1 13 12  DLIM 
DDG 14 15  DCGD 
R2 12 15 1 
D2 30 15  DLIM 
DSD 10 3  DSUB 
.MODEL PMOS PMOS  LEVEL = 3  U0 = 400  VMAX = 1E+006  ETA = 0.001 
+ TOX = 6E-008  NSUB = 1E+016  KP = 1.095  KAPPA = 49.86  VTO = -0.8823 
.MODEL DCGD D  CJO = 1.311E-011  VJ = 0.2302  M = 0.2576 
.MODEL DSUB D  IS = 3E-009  N = 1.688  RS = 0.5  BV = 25  CJO = 6.498E-012  VJ = 0.3007  M = 0.2934 
.MODEL DLIM D  IS = 0.0001 
.ENDS

*Diodes DMC2400UV Spice Model v1.0 Last Revised 2014/11/18