*---------- DMG3420U Spice Model ----------
.SUBCKT DMG3420U 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3  NMOS  L = 1E-006  W = 1E-006 
RD 10 1 0.02158 
RS 30 3 0.001 
RG 20 2 1.53 
CGS 2 3 3.785E-010 
EGD 12 0 2 1 1 
VFB 14 0 0 
FFB 2 1  VFB 1 
CGD 13 14 6.25E-010 
R1 13 0 1 
D1 12 13  DLIM 
DDG 15 14  DCGD 
R2 12 15 1 
D2 15 0  DLIM 
DSD 3 10  DSUB 
.MODEL NMOS NMOS  LEVEL = 3  VMAX = 1E+006  ETA = 0.009674  VTO = 1.32 
+ TOX = 6E-008  NSUB = 1E+016  KP = 53.82  KAPPA = 1E-015  U0 = 400 
.MODEL DCGD D  CJO = 3.069E-010  VJ = 0.1752  M = 0.4052 
.MODEL DSUB D  IS = 8.863E-010  N = 1.372  RS = 0.01813  BV = 22  CJO = 4.022E-011  VJ = 0.2305  M = 0.4418 
.MODEL DLIM D  IS = 0.0001 
.ENDS
*Diodes DMG3420U Spice Model v1.0 Last Revised 2010/5/9