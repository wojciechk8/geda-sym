*
*******************************************
*
*RB521S30
*
*NXP Semiconductors
*
*Schottky barrier rectifier
*
*
*
*
*IFSM = 1A    @ tp = 8,3ms
*VF   = 500mV @ IF = 0,2A
*
*
*
*
*
*
*
*
*
*
*Package pinning does not match Spice model pinning.
*Package: SOD523
*
*Package Pin 1: Cathode 
*Package Pin 2: Anode    
*     
*
*
*
*Simulator: SPICE3
*
*******************************************
*#
.SUBCKT RB521S30 1 2
*
* The resistor does not 
* reflect a physical device. 
* Instead it improves modeling
* in the reverse mode of 
* operation.
*
R1 1 2 4.771E+06
D1 1 2 RB521S30
*
.MODEL RB521S30 D
+ IS = 9.539E-07
+ N = 1.007
+ BV = 35
+ IBV = 0.001
+ RS = 0.4678
+ CJO = 3.518E-11
+ VJ = 0.3193
+ M = 0.4687
+ FC = 0.5
+ EG = 0.69
+ XTI = 2
.ENDS
*

