* TLC27L2 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.03 ON 07/10/90 AT 15:01
* REV (N/A)      SUPPLY VOLTAGE: 5V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TLC27L2  1 2 3 4 5
*
  C1   11 12 10.12E-12
  C2    6  7 15.00E-12
  CPSR 85 86 79.6E-9
  DCM+ 81 82 DX
  DCM- 83 81 DX
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  ECMR 84 99 (2,99)  1
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  EPSR 85 0 POLY(1) (3,4) -8.5E-6  1.7E-6
  ENSE 89 2 POLY(1) (88,0) 170E-6  1
  FB 7 99 POLY(6) VB VC VE VLP VLN VPSR 0 419.1E6 -70E6 70E6 70E6 -70E6 492E6
  GA    6  0 11 12 7.069E-6
  GCM 0  6 10 99 282.0E-12
  GPSR 85 86 (85,86) 100E-6
  GRD1 60 11 (60,11) 7.067E-6
  GRD2 60 12 (60,12) 7.067E-6
  HLIM 90  0 VLIM 1K
  HCMR 80 1 POLY(2) VCM+ VCM- 0 1E2 1E2
  IRP 3 4 9.55E-6
  ISS   3 10 DC 450.0E-9
  IIO 2 0 .1E-12
  I1 88 0 1E-21
  J1   11  89 10 JX
  J2   12  80 10 JX
  R2    6  9 100.0E3
  RCM 84 81 1K
  RN1 88 0 195E3
  RO1   8  5 85
  RO2   7 99 85
  RSS  10 99 444.4E6
  VAD  60 4 -.4
  VCM+ 82 99 1.1
  VCM- 83 99 -2.3
  VB    9  0 DC 0
  VC 3 53 DC 1.470
  VE   54  4 DC .57
  VLIM  7  8 DC 0
  VLP  91  0 DC 20
  VLN   0 92 DC 20
  VPSR 0 86 DC 0
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=300.0E-15 BETA=222.1E-6 VTO=.026 KF=1.45E-17)
.ENDS
