***** NE5532 Source: Texas Instruments NE5534
* C2 added to simulate compensated frequency response (Uwe Beis)

* NE5532 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING NE5534 model from Texas InstrumentsAT 12:41
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT NE5532   1 2 3 4 5
*
  C1   11 12 7.703E-12
  C2    6  7 23.500E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  FB    7 99 POLY(5) VB VC VE VLP VLN 0 2.893E6 -3E6 3E6 3E6 -3E6
  GA    6  0 11 12 1.382E-3
  GCM   0  6 10 99 13.82E-9
  IEE  10  4 DC 133.0E-6
  HLIM 90  0 VLIM 1K
  Q1   11  2 13 QX
  Q2   12  1 14 QX
  R2    6  9 100.0E3
  RC1   3 11 723.3
  RC2   3 12 723.3
  RE1  13 10 329
  RE2  14 10 329
  REE  10 99 1.504E6
  RO1   8  5 50
  RO2   7 99 25
  RP    3  4 7.757E3
  VB    9  0 DC 0
  VC    3 53 DC 2.700
  VE   54  4 DC 2.700
  VLIM  7  8 DC 0
  VLP  91  0 DC 38
  VLN   0 92 DC 38
.MODEL DX D(IS=800.0E-18)
.MODEL QX NPN(IS=800.0E-18 BF=132)
.ENDS
