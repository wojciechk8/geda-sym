.SUBCKT BSD840N_L0  drain  gate  source

Lg     gate  g1    1n
Ld     drain d1    0.5n
Ls     source s1   1n
Rs      s1    s2   46.66m

Rg     g1    g2     10.5
M1      d2    g2    s2    s2    DMOS    L=1u   W=1u
.MODEL DMOS NMOS ( KP= 7.5  VTO=1.17  THETA=0  VMAX=1.5e5  ETA=0.003  LEVEL=3)
Rd     d1    d2    121.71m TC=6.5m

Dbd     s2    d2    Dbt
.MODEL     Dbt    D(BV=24   M=0.35  CJO=0.03n  VJ=0.7V)
Dbody   s2   21    DBODY
.MODEL DBODY  D(IS=9.6p  N=1.21  RS=120.75u  EG=1.12  TT=3n)
Rdiode  d1  21    120.75m TC=7m

.MODEL   sw    NMOS(VTO=0  KP=10   LEVEL=1)
Maux      g2   c    a    a   sw
Maux2     b    d    g2    g2   sw
Eaux      c    a    d2    g2   1
Eaux2     d    g2   d2    g2   -1
Cox       b    d2   0.04n
.MODEL     DGD    D(M=1.1   CJO=0.04n   VJ=0.5)
Rpar      b    d2   1Meg
Dgd       a    d2   DGD
Rpar2     d2   a    10Meg
Cgs     g2    s2    0.05n

.ENDS  BSD840N_L0
